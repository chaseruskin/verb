import godan::*;

interface add_bfm #(
    parameter integer WORD_SIZE = 17
);
    logic cin;
    logic[WORD_SIZE-1:0] in0;
    logic[WORD_SIZE-1:0] in1;
    logic[WORD_SIZE-1:0] sum;
    logic cout;
endinterface

module add_tb #(
    parameter integer WORD_SIZE = 17
);

    add_bfm #(.WORD_SIZE(WORD_SIZE)) bfm();
    add_bfm #(.WORD_SIZE(WORD_SIZE)) mdl();

    add #(
        .WORD_SIZE(WORD_SIZE)
    ) dut (
        .cin(bfm.cin),
        .in0(bfm.in0),
        .in1(bfm.in1),
        .sum(bfm.sum),
        .cout(bfm.cout)
    );

    int events = $fopen("events.log", "w");

    logic clk, halt;
    time period = 10;

    always begin
        spin_clock(clk, period, halt);
    end

    // This task is automatically @generated by Verb.
    // It is not intended for manual editing.
    task send(int fd);
        automatic string row = "";
        if(!$feof(fd)) begin
            $fgets(row, fd);

            $sscanf(drive(row), "%b", bfm.cin);
            $sscanf(drive(row), "%b", bfm.in0);
            $sscanf(drive(row), "%b", bfm.in1);
        end
    endtask

    always begin: producer 
        int inputs = $fopen("inputs.txt", "r");
        while(!$feof(inputs)) begin
            send(inputs);
            @(posedge clk);
        end
        $fclose(inputs);
        wait(0);
    end

    // This task is automatically @generated by Verb.
    // It is not intended for manual editing.
    task compare(int fd);
        string row, rec, exp;
        if(!$feof(fd)) begin
            $fgets(row, fd);

            $sscanf(load(row), "%b", mdl.sum);
            $sformat(rec, "%b", bfm.sum);
            $sformat(exp, "%b", mdl.sum);
            assert_eq(events, rec, exp, "sum");

            $sscanf(load(row), "%b", mdl.cout);
            $sformat(rec, "%b", bfm.cout);
            $sformat(exp, "%b", mdl.cout);
            assert_eq(events, rec, exp, "cout");
        end
    endtask;

    always begin: consumer
        int outputs = $fopen("outputs.txt", "r");
        while(!$feof(outputs)) begin
            @(posedge clk);
            compare(outputs);
        end
        $fclose(outputs);
        complete(halt, events);
    end

endmodule