-- Project: Vertex
-- Package: tutils
--
-- Provides test utility functions for testbench simulation. This involves
-- reading interface signals, loading expected values, and various 
-- simulation-specific tasks.

library ieee;
use ieee.std_logic_1164.all;

library amp;
use amp.types.all;
use amp.cast.all;

library std;
use std.textio.all;

package tutils is

  -- Generates a half duty cycle clock `clk` with a period of `period` that
  -- is continuously driven until `halt` is set to true. 
  procedure spin_clock(signal clk: out logic; period: time; signal halt: bool);

  -- Asynchronously triggers the reset (active-high) and then synchronously
  -- deactivates the reset after `cycles` clock cycles generated by `clk`.
  --
  -- The reset will not be applied if `cycles` is set to 0. The reset will
  -- deactivate on the falling edge of the `cycles` count clock cycle.
  procedure trigger_reset_h(signal clk: logic; signal rst: out logic; cycles: usize);

  -- Asynchronously triggers the reset (active-low) and then synchronously
  -- deactivates the reset after `cycles` clock cycles generated by `clk`.
  --
  -- The reset will not be applied if `cycles` is set to 0. The reset will
  -- deactivate on the falling edge of the `cycles` count clock cycle.
  procedure trigger_reset_l(signal clk: logic; signal rst: out logic; cycles: usize);

  -- Drive a logic vector signal `x` with a value from the line `row`.
  procedure drive(variable row: inout line; signal x: out logics);

  -- Drive a logic bit signal `x` with a value from the line `row`.
  procedure drive(variable row: inout line; signal x: out logic);

  -- Read a logic vector value from the line `row` into the variable `x`.
  procedure load(variable row: inout line; variable x: out logics);

  -- Read a logic bit value from the line `row` into the variable `x`.
  procedure load(variable row: inout line; variable x: out logic);
  
  -- Sets `halt` to true and enters an infinite wait statement to signal 
  -- that the simulation is complete.
  procedure complete(signal halt: out bool);

  -- Enters an infinite wait if the `halt` signal is set to true.
  procedure check(halt: in bool);

  -- Awaits the flag to be asserted or until delay time is up. Sets `timeout`
  -- to true when the flag was asserted before the timeout and false if
  -- the timeout was reached before the flag was raised.
  --
  -- Sets an unbounded waiting limit if `cycles` is set to 0.
  procedure monitor_h(signal clk: logic; signal flag: logic; cycles: usize; variable timeout: out bool);

end package;


package body tutils is

  procedure complete(signal halt: out bool) is
  begin
    halt <= true;
    wait;
  end procedure;


  procedure check(halt: in bool) is
  begin
    if halt = true then 
      wait;
    end if;
  end procedure;


  procedure spin_clock(signal clk: out logic; period: time; signal halt: bool) is
    variable inner_clk : logic := '0';
  begin
    while halt = false loop
      clk <= inner_clk;
      wait for period/2;
      inner_clk := not inner_clk;
    end loop;
    wait;
  end procedure;


  procedure trigger_reset_h(signal clk: logic; signal rst: out logic; cycles: usize) is
  begin
    -- only apply the reset if the number of cycles to delay is greater than zero
    if cycles > 0 then
      rst <= '1';
      wait for 0 ns;
      for delay in 1 to cycles loop
        wait until rising_edge(clk);
      end loop;
      wait until falling_edge(clk);
    end if;
    rst <= '0';
    -- wait for 0 ns;
  end procedure;


  procedure trigger_reset_l(signal clk: logic; signal rst: out logic; cycles: usize) is
  begin
    -- only apply the reset if the number of cycles to delay is greater than zero
    if cycles > 0 then
      rst <= '0';
      wait for 0 ns;
      for delay in 1 to cycles loop
        wait until rising_edge(clk);
      end loop;
      wait until falling_edge(clk);
    end if;
    rst <= '1';
    -- wait for 0 ns;
  end procedure;


  procedure monitor_h(signal clk: logic; signal flag: logic; cycles: usize; variable timeout: out bool) is
    variable cycle_count : usize := 0;
  begin
    timeout := true;
    if cycles = 0 then
      wait until rising_edge(clk) and flag = '1';
      timeout := false;
    else
      while cycle_count < cycles loop
        if flag = '1' then
          timeout := false;
          exit;
        end if;
        wait until rising_edge(clk);
        cycle_count := cycle_count + 1;
      end loop;
    end if;
  end procedure;


  procedure drive(variable row: inout line; signal x: out logics) is
    variable word: str(x'range);
    variable temp: logics(x'range);
    variable delim: char;
  begin
    if row'length > 0 then
      read(row, word);
      for i in x'range loop
        temp(i) := to_logic(word(i));
      end loop;
      x <= temp;
      -- ignore the delimiter
      read(row, delim);
      -- wait for 0 ns;
    end if;
  end procedure;


  procedure load(variable row: inout line; variable x: out logics) is
    variable word: str(x'range);
    variable delim: char;
  begin
    if row'length > 0 then
      read(row, word);
      for i in x'range loop
        x(i) := to_logic(word(i));
      end loop;
      -- ignore the delimiter
      read(row, delim);
    end if;
  end procedure;


  procedure drive(variable row: inout line; signal x: out logic) is
    variable word: char;
    variable delim: char;
  begin
    if row'length > 0 then
      read(row, word);
      x <= to_logic(word);
      -- ignore the delimiter
      read(row, delim);
      -- wait for 0 ns;
    end if;
  end procedure;


  procedure load(variable row: inout line; variable x: out logic) is
      variable word: char;
      variable delim: char;
  begin
    if row'length > 0 then
      read(row, word);
      x := to_logic(word);
      -- ignore the delimiter
      read(row, delim);
    end if;
  end procedure;

end package body;